/*---------------------------------------------------------------------------
 *
 *  Copyright (c) 2023 by Jin Hyeong Park, All rights reserved.
 *
 *  File name  : Fadder_Fsubtractor.v
 *  Written by : Park, Jin Hyoeng
 *               School of Electrical Engineering / Department of Biomechatronics
 *               Sungkyunkwan University
 *  Written on : January 18, 2023
 *  Version    : 2.0
 *  Design     : Floating Point Number Adder and Subtractor
 *  Target Devices: Zybo Z7-20
 *  Modification History:
 *      * January 10, 2023  Jin Hyeong Park
 *        version 1.0 released.
 *
 *      * January 18, 2023 by Jin Hyeong Park
 *        version 2.0 released.
 *
 *      * January 25, 2023 by Jin Hyeong Park
 *        version 2.0 code modified and comments added.
 *
 *  NOTE: Overflow and Underflow are not considered yet.
 *
 *---------------------------------------------------------------------------*/


module Fadder_Fsubtractor(
    input clk,
    input [31:0] A,
    input [31:0] B,
    input reset_n,
    output reg [31:0] result
);

reg result_sign;
reg [7:0] result_exponent;
reg [22:0] result_fraction;

// A and B - sign, exponent, fraction 
reg A_sign, B_sign;
reg [7:0] A_exponent, B_exponent;
reg [22:0] A_fraction, B_fraction;

// Big and Small - sign, exponent, fraction
reg big_sign, small_sign;
reg [7:0] big_exponent, small_exponent;
reg [22:0] big_fraction, small_fraction;

// Difference
reg [7:0] exponent_diff;
reg input_diff;

// Temp Big Fraction & Temp Small Fraction & Temp Fraction
reg [23:0] tb_fraction, ts_fraction, temp_fraction;
// Temp Exponent
reg [7:0] temp_exponent;
reg carry;

always @ (posedge clk) begin
    A_sign = A[31];
    B_sign = B[31];
    A_exponent = A[30:23];
    B_exponent = B[30:23];
    A_fraction = A[22:0];
    B_fraction = B[22:0];
    
    input_diff = ({A_exponent, A_fraction} >= {B_exponent, B_fraction}) ? 1'b1 : 1'b0;
    exponent_diff = A_exponent - B_exponent;
    big_sign = (input_diff) ? A_sign : B_sign;
    big_exponent = (input_diff) ? A_exponent : B_exponent;
    big_fraction = (input_diff) ? A_fraction : B_fraction;
    
    small_sign = (input_diff) ? B_sign : A_sign;
    small_exponent = (input_diff) ? B_exponent : A_exponent;
    small_fraction = (input_diff) ? B_fraction : A_fraction;
    
    tb_fraction = {1'b1, big_fraction};
    ts_fraction = {1'b1, small_fraction};
    ts_fraction = ts_fraction >> exponent_diff;
    
    {carry, temp_fraction} = (big_sign == small_sign) ? tb_fraction + ts_fraction : tb_fraction - ts_fraction;

    temp_exponent = big_exponent;
    
    if (!reset_n) begin
        temp_fraction = 0;
        temp_exponent = 0;
    end else begin
        if (carry) begin
            temp_fraction = temp_fraction >> 1'b1;
            temp_exponent = temp_exponent + 1'b1;
        end else begin
            if (!temp_fraction[23]) begin
                temp_fraction = temp_fraction << 1;
                temp_exponent = temp_exponent - 1'b1;
            end else begin
                temp_fraction = temp_fraction;
                temp_exponent = temp_exponent;
            end
        end
    end

    result_sign = big_sign;
    result_fraction = temp_fraction[22:0];
    result_exponent = temp_exponent;
    result = {result_sign, result_exponent, result_fraction};
end

endmodule
