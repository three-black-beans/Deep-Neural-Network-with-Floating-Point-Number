module DNN_tb();

reg clk = 0;
reg [31:0] x1, x2, x3;
reg set;
reg [31:0] target_out;

wire [31:0] out;
wire [2:0] control;

neural_network tb(.control(control), .target_out(target_out), .clk(clk), .x1(x1), .x2(x2), .x3(x3), .out(out), .set(set));

always #1
clk = ~clk;

initial begin
    x1 = 0;
    x2 = 0;
    x3 = 0;
    target_out = 0;
    set = 1;
    
    #11
    set = 0;

    repeat(500000) begin
    #12

    x1 = 32'b00111111100000000000000000000000;
    x2 = 32'b00111111100000000000000000000000;
    x3 = 32'b00111111100000000000000000000000;
    target_out = 32'b00111111010000000000000000000000;

    #12
    x1 = 32'b01000000010000000000000000000000;
    x2 = 32'b01000000010000000000000000000000;
    x3 = 32'b01000000010000000000000000000000;
    target_out = 32'b00111111000000000000000000000000;

    #12
    x1 = 32'b01000000110000000000000000000000;
    x2 = 32'b01000000110000000000000000000000;
    x3 = 32'b01000000110000000000000000000000;
    target_out = 32'b00111110110000000000000000000000;
    
    end
end

endmodule